-- Genereert een sinus van ~1KHz (of gespecificeerde 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY toongenerator IS
	GENERIC (wait_cycles : natural := 800);

	PORT(
		clock, activate : IN std_logic;
		data : OUT std_logic_vector(15 downto 0)
	);
END toongenerator;

ARCHITECTURE behaviour OF toongenerator IS
	FUNCTION sinlut (n:std_logic_vector(5 DOWNTO 0)) RETURN std_logic_vector IS BEGIN
		CASE n IS  -- 6 bits to 2s complement 16 bit sine wave
			WHEN "000000" => RETURN "0000000000000000";
			WHEN "000001" => RETURN "0000001100100010";
			WHEN "000010" => RETURN "0000011000111101";
			WHEN "000011" => RETURN "0000100101001000";
			WHEN "000100" => RETURN "0000110000111101";
			WHEN "000101" => RETURN "0000111100010011";
			WHEN "000110" => RETURN "0001000111000101";
			WHEN "000111" => RETURN "0001010001001010";
			WHEN "001000" => RETURN "0001011010011110";
			WHEN "001001" => RETURN "0001100010111001";
			WHEN "001010" => RETURN "0001101010011000";
			WHEN "001011" => RETURN "0001110000110110";
			WHEN "001100" => RETURN "0001110110001110";
			WHEN "001101" => RETURN "0001111010011101";
			WHEN "001110" => RETURN "0001111101100001";
			WHEN "001111" => RETURN "0001111111010111";
			WHEN "010000" => RETURN "0001111111111111";
			WHEN "010001" => RETURN "0001111111011000";
			WHEN "010010" => RETURN "0001111101100011";
			WHEN "010011" => RETURN "0001111010100001";
			WHEN "010100" => RETURN "0001110110010011";
			WHEN "010101" => RETURN "0001110000111100";
			WHEN "010110" => RETURN "0001101010100000";
			WHEN "010111" => RETURN "0001100011000010";
			WHEN "011000" => RETURN "0001011010100111";
			WHEN "011001" => RETURN "0001010001010100";
			WHEN "011010" => RETURN "0001000111001111";
			WHEN "011011" => RETURN "0000111100011111";
			WHEN "011100" => RETURN "0000110001001001";
			WHEN "011101" => RETURN "0000100101010101";
			WHEN "011110" => RETURN "0000011001001010";
			WHEN "011111" => RETURN "0000001100101111";
			WHEN "100000" => RETURN "0000000000001101";
			WHEN "100001" => RETURN "1111110011101010";
			WHEN "100010" => RETURN "1111100111010000";
			WHEN "100011" => RETURN "1111011011000100";
			WHEN "100100" => RETURN "1111001111001110";
			WHEN "100101" => RETURN "1111000011111000";
			WHEN "100110" => RETURN "1110111001000110";
			WHEN "100111" => RETURN "1110101111000000";
			WHEN "101000" => RETURN "1110100101101100";
			WHEN "101001" => RETURN "1110011101001110";
			WHEN "101010" => RETURN "1110010101101110";
			WHEN "101011" => RETURN "1110001111010000";
			WHEN "101100" => RETURN "1110001001110110";
			WHEN "101101" => RETURN "1110000101100110";
			WHEN "101110" => RETURN "1110000010100010";
			WHEN "101111" => RETURN "1110000000101010";
			WHEN "110000" => RETURN "1110000000000000";
			WHEN "110001" => RETURN "1110000000100110";
			WHEN "110010" => RETURN "1110000010011010";
			WHEN "110011" => RETURN "1110000101011010";
			WHEN "110100" => RETURN "1110001001101000";
			WHEN "110101" => RETURN "1110001110111110";
			WHEN "110110" => RETURN "1110010101011000";
			WHEN "110111" => RETURN "1110011100110110";
			WHEN "111000" => RETURN "1110100101010000";
			WHEN "111001" => RETURN "1110101110100010";
			WHEN "111010" => RETURN "1110111000100110";
			WHEN "111011" => RETURN "1111000011010110";
			WHEN "111100" => RETURN "1111001110101010";
			WHEN "111101" => RETURN "1111011010011110";
			WHEN "111110" => RETURN "1111100110101010";
			WHEN OTHERS   => RETURN "1111110011000100";
			END CASE;
	END sinlut;  

	SIGNAL index : unsigned(5 downto 0) := (OTHERS => '0');

BEGIN 
	PROCESS (clock, activate) 
		VARIABLE wait_counter : integer RANGE 0 TO wait_cycles := 0;
	BEGIN  
		IF rising_edge(clock) AND activate = '1' THEN
			IF wait_counter = wait_cycles THEN
				wait_counter <= 0;        
				index <= index + 1;
			ELSE
				wait_counter <= wait_counter + 1;
			END IF;
		END IF;
	END PROCESS;

	data <= sinlut(std_logic_vector(index));

END behaviour;